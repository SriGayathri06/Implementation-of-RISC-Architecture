`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:34:10 03/02/2022 
// Design Name: 
// Module Name:    pc_assign 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// File: pc_assign.v
// Generated by MyHDL 0.11
// Date: Wed Mar  2 16:10:07 2022


`timescale 1ns/10ps

module pc_assign (
    input reset,
    output reg [31:0] read_addr,
    input [31:0] pc
);

/*
input reset;
output [31:0] read_addr;
reg [31:0] read_addr;
input [31:0] pc;
*/



always @(*) begin: PC_ASSIGN_ASSIGN
    if ((reset == 1)) begin
        read_addr = pc;
    end
    //
    else 
        read_addr = 32'bX;
    //
end

endmodule

