`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:32:39 03/02/2022 
// Design Name: 
// Module Name:    alu_control 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// File: alu_control.v
// Generated by MyHDL 0.11
// Date: Wed Mar  2 16:10:07 2022


`timescale 1ns/10ps

module alu_control (
    reset,
    instruction,
    alu_op,
    alu_decode
);

input reset;
input [31:0] instruction;
input [3:0] alu_op;
output [3:0] alu_decode;
reg [3:0] alu_decode1;




always @(instruction,reset,alu_op) begin: ALU_CONTROL_ALUCONT
    if ((reset == 1)) begin
        case (alu_op)
            'h2: begin
                if ((instruction[32-1:25] == 0)) begin
                    if ((instruction[15-1:12] == 0)) begin
                        alu_decode1 <= 2;
                    end
                    else if ((instruction[15-1:12] == 1)) begin
                        alu_decode1 <= 3;
                    end
                    else if ((instruction[15-1:12] == 2)) begin
                        alu_decode1 <= 4;
                    end
                    else if ((instruction[15-1:12] == 3)) begin
                        alu_decode1 <= 5;
                    end
                    else if ((instruction[15-1:12] == 4)) begin
                        alu_decode1<=7;
                    end
                    else if ((instruction[15-1:12] == 5)) begin
                        alu_decode1 <= 8;
                    end
                    else if ((instruction[15-1:12] == 6)) begin
                        alu_decode1 <= 1;
                    end
                    else if ((instruction[15-1:12] == 7)) begin
                        alu_decode1 <= 0;
                    end
                    //
                    else
                        alu_decode1<=4'bX;
                    //
                end
                else if ((instruction[32-1:25] == 32)) begin
                    if ((instruction[15-1:12] == 0)) begin
                        alu_decode1 <= 6;
                    end
                    else if ((instruction[15-1:12] == 5)) begin
                        alu_decode1 <= 9;
                    end
                    else
                        alu_decode1<=4'bX;
                end
                //
                else
                    alu_decode1<=4'bx;
                //
            end
            'h0: begin
                alu_decode1 <= 2;
            end
            'h7: begin
                if ((instruction[15-1:12] == 0)) begin
                    alu_decode1 <= 7;
                end
                //
                else
                    alu_decode1<=4'bX;
                //
            end
            default: 
                alu_decode1<=4'bX;
        endcase
    end
    //
    else 
        alu_decode1<=4'bX;
    //
end
assign alu_decode=alu_decode1;
endmodule

