`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:33:26 03/02/2022 
// Design Name: 
// Module Name:    imm_gen 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// File: imm_gen.v
// Generated by MyHDL 0.11
// Date: Wed Mar  2 16:10:07 2022


`timescale 1ns/10ps

module imm_gen (
    reset,
    instruction,
    im_gen
);


input reset;
input [31:0] instruction;
output [31:0] im_gen;
reg [31:0] im_gen1;


reg [31:0]x;

always @(instruction, reset) begin: IMM_GEN_IMMGEN
    //integer temp;
    if ((reset == 1)) begin
        if ((instruction[7-1:0] == 3)) begin
            im_gen1[12-1:0] <= instruction[32-1:20];
        end
        else if ((instruction[7-1:0] == 35)) begin
            im_gen1[12-1:5] <= instruction[32-1:25];
            im_gen1[5-1:0] <= instruction[12-1:7];
        end
        else if ((instruction[7-1:0] == 99)) begin
            im_gen1[12] <= instruction[31];
            im_gen1[11-1:5] <= instruction[31-1:25];
            im_gen1[11] <= instruction[7];
            im_gen1[5-1:1] <= instruction[12-1:8];
            im_gen1[0] <= 0;
        end
        //
        else
            im_gen1<=32'bX;
        //
        if ((instruction[31] == 0)) begin
            x=32'd0;
            im_gen1[32-1:(31 - 20)+1] <= x[19:0];
        end
        else if ((instruction[31] == 1))  begin
            //temp = ((2 ** 20) - 1);
			x=32'd1048575;
            im_gen1[32-1:(31 - 20)+1] <= x[19:0];
        end
        else 
            im_gen1<=32'bX;
    end
    //
    else
        im_gen1<=32'bX;
    //
end
assign im_gen=im_gen1;
endmodule

