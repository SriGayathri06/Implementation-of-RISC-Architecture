`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:19:43 03/02/2022 
// Design Name: 
// Module Name:    control 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// File: control.v
// Generated by MyHDL 0.11
// Date: Wed Mar  2 16:10:06 2022


`timescale 1ns/10ps

module control (
    
    reset,
    opcode,
    brnch,
    mem_rd,
    mem_to_rgs,
    alu_op,
    mem_wr,
    alu_src,
    reg_wr
);


input reset;
input [6:0] opcode;
output [0:0] brnch;
reg [0:0] brnch1;
output [0:0] mem_rd;
reg [0:0] mem_rd1;
output [0:0] mem_to_rgs;
reg [0:0] mem_to_rgs1;
output [3:0] alu_op;
reg [3:0] alu_op1;
output [0:0] mem_wr;
reg [0:0] mem_wr1;
output [0:0] alu_src;
reg [0:0] alu_src1;
output [0:0] reg_wr;
reg [0:0] reg_wr1;




always @(opcode, reset) begin: CONTROL_CONT
    if ((reset == 1)) begin
        case (opcode)
            'h33: begin
                alu_src1 <= 1'b0;
                mem_to_rgs1 <= 1'b0;
                reg_wr1 <= 1'b1;
                mem_rd1 <= 1'b0;
                mem_wr1 <= 1'b0;
                brnch1 <= 1'b0;
                alu_op1 <= 2;
            end
            'h3: begin
                alu_src1 <= 1'b1;
                mem_to_rgs1 <= 1'b1;
                reg_wr1 <= 1'b1;
                mem_rd1 <= 1'b0;
                mem_wr1 <= 1'b0;
                brnch1 <= 1'b0;
                alu_op1 <= 0;
            end
            'h23: begin
                alu_src1 <= 1'b1;
                mem_to_rgs1 <= 1'b0;
                reg_wr1 <= 1'b0;
                mem_rd1 <= 1'b0;
                mem_wr1 <= 1'b1;
                brnch1 <= 1'b0;
                alu_op1 <= 0;
            end
            'h63: begin
                alu_src1 <= 1'b0;
                mem_to_rgs1 <= 1'b0;
                reg_wr1 <= 1'b0;
                mem_rd1 <= 1'b0;
                mem_wr1 <= 1'b0;
                brnch1 <= 1'b1;
                alu_op1 <= 7;
            end
            default:begin
                alu_src1 <= 1'bX;
                mem_to_rgs1 <= 1'bX;
                reg_wr1 <= 1'bX;
                mem_rd1 <= 1'bX;
                mem_wr1 <= 1'bX;
                brnch1<= 1'bX;
                alu_op1 <= 4'bX;
            end
            endcase
    end
    //
    else begin
        alu_src1 <= 1'bX;
        mem_to_rgs1 <= 1'bX;
        reg_wr1 <= 1'bX;
        mem_rd1 <= 1'bX;
        mem_wr1 <= 1'bX;
        brnch1 <= 1'bX;
        alu_op1 <= 4'bX;
    end
end
assign alu_src=alu_src1 ;
assign mem_to_rgs=mem_to_rgs1 ;
assign reg_wr=reg_wr1 ;
assign mem_rd=mem_rd1 ;
assign mem_wr=mem_wr1 ;
assign brnch=brnch1 ;
assign alu_op=alu_op1;

endmodule

