`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:32:00 03/02/2022 
// Design Name: 
// Module Name:    wda_mux 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// File: wda_mux.v
// Generated by MyHDL 0.11
// Date: Wed Mar  2 16:10:07 2022


`timescale 1ns/10ps

module wda_mux (
    reset,
    wda,
    mem_to_rgs,
    result,
    read_data
);


input reset;
output [31:0] wda;
reg [31:0] wda1;
input [0:0] mem_to_rgs;
input [31:0] result;
input [31:0] read_data;




always @(mem_to_rgs, reset,read_data,result) begin: WDA_MUX_WMUX
    if ((reset == 1)) begin
        if (mem_to_rgs) begin
            wda1 <= read_data;
        end
        else begin
            wda1 <= result;
        end
    end
    //
    else
        wda1=32'dX;
    //
end
assign wda=wda1;
endmodule

