`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:29:50 03/02/2022 
// Design Name: 
// Module Name:    alu_mux 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// File: alu_mux.v
// Generated by MyHDL 0.11
// Date: Wed Mar  2 16:10:07 2022


`timescale 1ns/10ps

module alu_mux (
    reset,
    im_gen,
    rdb,
    rdx,
    alu_src
);


input reset;
input [31:0] im_gen;
input [31:0] rdb;
output [31:0] rdx;
reg [31:0] rdx1;
input [0:0] alu_src;




always @(reset,im_gen,rdb,alu_src) begin: ALU_MUX_AMUX
    if ((reset == 1)) begin
        if (alu_src) begin
            rdx1 <= im_gen;
        end
        else begin
            rdx1 <= rdb;
        end
    end
    //
    else
        rdx1<=32'bX;
    //
end
assign rdx=rdx1;
endmodule

