`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:34:45 03/02/2022 
// Design Name: 
// Module Name:    taken 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
// File: taken.v
// Generated by MyHDL 0.11
// Date: Wed Mar  2 16:10:07 2022


`timescale 1ns/10ps



module taken (
    result,
    brnch,
    pc_sel
);


input [31:0] result;
input [0:0] brnch;
output [0:0] pc_sel;
reg [0:0] pc_sel1;




always @(brnch, result) begin: TAKEN_TAKE
    if (((result == 0) & brnch)) begin
        pc_sel1 <= 1'b1;
    end
    else begin
        pc_sel1 <= 1'b0;
    end
end
assign pc_sel=pc_sel1;
endmodule

